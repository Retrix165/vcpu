module CPU(i_clk);

    input wire i_clk;

    parameter filepath = "";
    parameter numInstructions = 0;

    initial begin

    end

    always @(posedge i_clk) begin //datapath here probably
    
    end

endmodule